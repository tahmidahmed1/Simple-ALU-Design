-- ECE 124, LAB Session #206, Team Number #9, Tahmid Ahmed & Vidhi Patel
library ieee;
use ieee.std_logic_1164.all;

entity hex_mux is 
port ( 
	hex_num3, hex_num2, hex_num1, hex_num0 : in std_logic_vector(3 downto 0); -- 4-bit inputs
	mux_select										: in std_logic_vector(1 downto 0); -- 2-bit selector
	hex_out											: out std_logic_vector(3 downto 0) -- The hex output
);

end hex_mux;

architecture mux_logic of hex_mux is 

begin 

	-- for the multiplexing of four hex input busses 
	with mux_select(1 downto 0) select
	hex_out <= hex_num0 when "00", -- when input from mux_select is "00" hex_num0 will be selected.
				  hex_num1 when "01", -- when input from mux_select is "01" hex_num1 will be selected.
				  hex_num2 when "10", -- when input from mux_select is "10" hex_num2 will be selected.
				  hex_num3 when "11"; -- when input from mux_select is "11" hex_num3 will be selected.
				  
end mux_logic;
